

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO SYS_TOP 
  PIN SI[3] 
    ANTENNAPARTIALMETALAREA 0.269 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.29389 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.026 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.93746 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 11.948 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 57.6623 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 25.314 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 121.953 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 496.391 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 2401.43 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA56 ;
  END SI[3]
  PIN SI[2] 
    ANTENNAPARTIALMETALAREA 0.187 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.89947 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 11.829 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.0899 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 9.16 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 44.252 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 189.881 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 930.724 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA56 ;
  END SI[2]
  PIN SI[1] 
    ANTENNAPARTIALMETALAREA 0.341 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.64021 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.04906 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 18.976 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 91.6594 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 495.891 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 2402.45 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA56 ;
  END SI[1]
  PIN SI[0] 
    ANTENNAPARTIALMETALAREA 0.997 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.98797 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 21.3255 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 105.534 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.677298 LAYER VIA23 ;
  END SI[0]
  PIN SO[3] 
    ANTENNAPARTIALMETALAREA 0.199 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.95719 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 5.973 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 28.9225 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 1.737 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 16.458 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 79.3554 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0702 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 286.547 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 1303.78 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.05698 LAYER VIA56 ;
  END SO[3]
  PIN SO[2] 
    ANTENNADIFFAREA 1.431 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 1.342 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.45502 LAYER METAL3 ;
  END SO[2]
  PIN SO[1] 
    ANTENNAPARTIALMETALAREA 5.722 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.9076 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4108 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 40.565 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 196.241 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.351509 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL4 ;
    ANTENNAGATEAREA 0.4108 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 40.918 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 198.407 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 0.439387 LAYER VIA45 ;
    ANTENNADIFFAREA 1.737 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 26.602 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 128.34 LAYER METAL5 ;
    ANTENNAGATEAREA 0.4108 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 105.675 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 510.823 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.439387 LAYER VIA56 ;
  END SO[1]
  PIN SO[0] 
    ANTENNAPARTIALMETALAREA 0.199 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.95719 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 2.207 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.8081 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 1.737 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 30.644 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 147.59 LAYER METAL5 ;
  END SO[0]
  PIN scan_clk 
    ANTENNAPARTIALMETALAREA 0.337 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.62097 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.288 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.38768 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 0.55557 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 2.75522 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.0235732 LAYER VIA34 ;
  END scan_clk
  PIN scan_rst 
    ANTENNAPARTIALMETALAREA 0.305 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.46705 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 12.884 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 62.5492 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1066 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 163.433 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 791.673 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 2.37054 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.502 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 17.037 LAYER METAL4 ;
    ANTENNAGATEAREA 0.1599 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 185.335 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 898.221 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.37054 LAYER VIA45 ;
  END scan_rst
  PIN test_mode 
    ANTENNAPARTIALMETALAREA 0.287 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.38047 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.452 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.17652 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 23.4948 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 116.424 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.828932 LAYER VIA34 ;
  END test_mode
  PIN SE 
    ANTENNAPARTIALMETALAREA 0.237 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.13997 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.354 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.5151 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1755 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 19.2456 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 93.9882 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.411396 LAYER VIA34 ;
  END SE
  PIN RST_N 
    ANTENNAPARTIALMETALAREA 0.565 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.71765 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.206 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.99326 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 2.19 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7263 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 52.5328 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 260.046 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.03189 LAYER VIA45 ;
  END RST_N
  PIN UART_CLK 
    ANTENNAPARTIALMETALAREA 0.269 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.29389 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.714 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.62674 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.616 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.96536 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 1.08319 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 5.3559 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.0353598 LAYER VIA45 ;
  END UART_CLK
  PIN REF_CLK 
    ANTENNAPARTIALMETALAREA 0.373 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.79413 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.7542 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 0.716207 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 3.52789 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.0235732 LAYER VIA34 ;
  END REF_CLK
  PIN UART_RX_IN 
    ANTENNAPARTIALMETALAREA 0.341 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.64021 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.55 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8379 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 9.734 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 47.0129 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4693 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 99.0105 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 477.187 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.86304 LAYER VIA56 ;
  END UART_RX_IN
  PIN UART_TX_O 
    ANTENNADIFFAREA 1.737 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.736 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.1602 LAYER METAL3 ;
  END UART_TX_O
  PIN parity_error 
    ANTENNAPARTIALMETALAREA 0.85 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0885 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 5.823 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 28.201 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 1.737 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 25.15 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 121.164 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1833 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 217.882 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 1057.27 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.42578 LAYER VIA56 ;
  END parity_error
  PIN framing_error 
    ANTENNAPARTIALMETALAREA 0.199 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.95719 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.659 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.17219 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 1.737 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 29.332 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 141.279 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1833 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 250.659 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 1216.19 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.64635 LAYER VIA56 ;
  END framing_error
END SYS_TOP

END LIBRARY
